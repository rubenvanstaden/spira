* Inductances

* Ports
.end